module test();
int a,b;
initial
begin
	$display("the value of a %d and b %0d",a,b);
// new line is added
//new line addded
//this is V3
end
endmodule
