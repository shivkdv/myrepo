module test();
int a,b;
initial
begin
	$display("the value of a %d and b %0d",a,b);
end
endmodule
