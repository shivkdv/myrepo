module test();
  initial
    begin
      $display("this code is going to pull to local from remote");
    end
endmodule
