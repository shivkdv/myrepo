fnffnfsdfbsdjsdjfsd
